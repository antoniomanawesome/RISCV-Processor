//made alu package so it's easier to see what does what in alu.sv
package alu_pkg;
    typedef enum logic [5:0] {
        add   = 6'd0,
        sub   = 6'd1,
        sll   = 6'd2,
        srl   = 6'd3,
        sra   = 6'd4,
        aand  = 6'd5,
        oor    = 6'd6,
        xxor  = 6'd7,
        slt   = 6'd8,
        sltu  = 6'd9,
        addi  = 6'd10,
        slli  = 6'd11,
        srli  = 6'd12,
        srai  = 6'd13,
        andi  = 6'd14,
        ori   = 6'd15,
        xori  = 6'd16,
        slti  = 6'd17,
        sltiu = 6'd18,
        lui   = 6'd19,
        auipc = 6'd20,
        lb = 6'd21,
        lbu = 6'd22,
        lh = 6'd23,
        lhu = 6'd24,
        lw = 6'd25,
        sb = 6'd26,
        sh = 6'd27,
        sw = 6'd28,
        fence = 6'd29,
        fence_i = 6'd30,
        jal = 6'd31,
        jalr = 6'd32,
        beq = 6'd33,
        bne = 6'd34,
        blt = 6'd35,
        bge = 6'd36,
        bltu = 6'd37,
        bgeu = 6'd38
    } alu_sel_t;
endpackage