module controller_tb
(
    
);
endmodule