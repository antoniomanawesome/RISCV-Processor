//creating instruction memory (where we put our file with the things we want to run)

module imem
#(parameter int WIDTH = 32)
(
    input logic [WIDTH-1:0] addr, //byte address from the program counter
);

endmodule