module alu


endmodule