package alu_pkg;
    typedef enum logic [4:0] {
        add   = 5'd0,
        sub   = 5'd1,
        sll   = 5'd2,
        srl   = 5'd3,
        sra   = 5'd4,
        and   = 5'd5,
        or    = 5'd6,
        xor   = 5'd7,
        slt   = 5'd8,
        sltu  = 5'd9,
        addi  = 5'd10,
        slli  = 5'd11,
        srli  = 5'd12,
        srai  = 5'd13,
        andi  = 5'd14,
        ori   = 5'd15,
        xori  = 5'd16,
        slti  = 5'd17,
        sltiu = 5'd18,
        lui   = 5'd19,
        auipc = 5'd20,
    } alu_sel_t;
endpackage